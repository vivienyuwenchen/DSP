//-----------------------------------------------------------------------------
// Multiplier
//-----------------------------------------------------------------------------

module multiplier #( parameter W = 16 )
(
    input  [W-1:0]   a,
    input  [W-1:0]   b,
    output [W*2-1:0] out
);

	assign out = a * b;

endmodule
