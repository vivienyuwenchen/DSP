//-----------------------------------------------------------------------------
// Multiplexers
//-----------------------------------------------------------------------------

// Two-input MUX with parameterized bit width (default: 32-bits)
module mux2 #( parameter W = 32 )
(
    input[W-1:0]    in0,
    input[W-1:0]    in1,
    input           sel,
    output[W-1:0]   out
);

    // Conditional operator - http://www.verilog.renerta.com/source/vrg00010.htm
    assign out = (sel) ? in1 : in0;

endmodule

// Four-input MUX with parameterized bit width (default: 32-bits)
module mux4 #( parameter W = 32 )
(
    input [W-1:0] in0,              // 4-bit input called a
    input [W-1:0] in1,              // 4-bit input called b
    input [W-1:0] in2,              // 4-bit input called c
    input [W-1:0] in3,              // 4-bit input called d
    input [1:0] sel,                // input sel used to select between a,b,c,d
    output [W-1:0] out              // 4-bit output based on input sel
);

    // When sel[1] is 0, (sel[0]? b:a) is selected and when sel[1] is 1, (sel[0] ? d:c) is taken
    // When sel[0] is 0, a is sent to output, else b and when sel[0] is 0, c is sent to output, else d
    assign out = sel[1] ? (sel[0] ? in3 : in2) : (sel[0] ? in1 : in0);

endmodule

// Eight-input MUX with parameterized bit width (default: 32-bits)
module mux8 #( parameter W = 32 )
(
    input [W-1:0] in0, in1, in2, in3, in4, in5, in6, in7,
    input [2:0] sel,    
    output [W-1:0] out
);

    // When sel[2] is 0, (sel[1] ? d:c:b:a) is selected and when sel[2] is 1, (sel[1] ? h:g:f:e) is taken
    // When sel[1] is 0, (sel[0] ? b:a) is selected and when sel[1] is 1, (sel[0] ? d:c) is taken
    // When sel[0] is 0, a is sent to output, else b and when sel[0] is 0, c is sent to output, else d
    assign out = sel[2] ? (sel[1] ? (sel[0] ? in7 : in6) : (sel[0] ? in5 : in4)) : (sel[1] ? (sel[0] ? in3 : in2) : (sel[0] ? in1 : in0));

endmodule
